
--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   14:57:52 01/13/2016
-- Design Name:   
-- Module Name:   /home/csmajs/kchan049/lab1/tb.vhd
-- Project Name:  lab1
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: my_alu
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY tb IS
END tb;
 
ARCHITECTURE behavior OF tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT my_alu
    PORT(
         A : IN  std_logic_vector(7 downto 0);
         B : IN  std_logic_vector(7 downto 0);
         opcode : IN  std_logic_vector(2 downto 0);
         result : OUT  std_logic_vector(7 downto 0);
         carryout : OUT  std_logic;
         overflow : OUT  std_logic;
         zero : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal A : std_logic_vector(7 downto 0) := (others => '0');
   signal B : std_logic_vector(7 downto 0) := (others => '0');
   signal opcode : std_logic_vector(2 downto 0) := (others => '0');

 	--Outputs
   signal result : std_logic_vector(7 downto 0);
   signal carryout : std_logic;
   signal overflow : std_logic;
   signal zero : std_logic;
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: my_alu PORT MAP (
          A => A,
          B => B,
          opcode => opcode,
          result => result,
          carryout => carryout,
          overflow => overflow,
          zero => zero
        );

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
		-- unsigned add
		opcode <= "000";
		A <= "00000000";
		B <= "00000000";
		
		wait for 100 ns;
		
		opcode <= "000";
		A <= "11000100";
		B <= "00000000";
		
		wait for 100 ns;
		
		--- signed add
		opcode <= "001";
		A <= "00000000";
		B <= "00000000";
		
		wait for 100 ns;
		
		opcode <= "001";
		A <= "01000100";
		B <= "01000000";
		
		wait for 100 ns;
		
		opcode <= "001";
		A <= "11000100";
		B <= "01000000";
		
		wait for 100 ns;
		
		--unsigned sub
		
		opcode <= "010";
		A <= "01000100";
		B <= "01000000";
		
		wait for 100 ns;
		
		opcode <= "010";
		A <= "00000100";
		B <= "01000000";
		
		wait for 100 ns;
		
		--signed sub
		
		opcode <= "011";
		A <= "01000100";
		B <= "01000000";
		
		
		wait for 100 ns;
		
		opcode <= "011";
		A <= "00000100";
		B <= "00000100";
		
		wait for 100 ns;
		
		opcode <= "011";
		A <= "00000100";
		B <= "01000000";
		
		wait for 100 ns;
		
		--and
		
		opcode <= "100";
		A <= "01000100";
		B <= "01000000";
		
		wait for 100 ns;
		
		opcode <= "100";
		A <= "00000100";
		B <= "01000000";
		
		wait for 100 ns;
		
		--or
		
		opcode <= "100";
		A <= "01000100";
		B <= "01000000";
		
		wait for 100 ns;
		
		opcode <= "100";
		A <= "00000000";
		B <= "00000000";
		
		wait for 100 ns;
		
		--xor
		
		opcode <= "110";
		A <= "01000100";
		B <= "01000000";
		
		wait for 100 ns;
		
		opcode <= "110";
		A <= "00000000";
		B <= "00000000";
		
		wait for 100 ns;
		
		--divide by 2
		opcode <= "111";
		A <= "00000100";
		
		wait for 100 ns;
		
		opcode <= "111";
		A <= "11000100";
		
		wait for 100 ns;

      wait;
   end process;

END;
